package sfifo_sequence_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	import sfifo_agent_pkg::*;
	`include "sfifo_sequence.svh"
endpackage